0.4 0.4 0.9 
0.2 0.2 0.2 
0.5 0.5 0.5 
1 1 1 
0.05 0.05 0.05 
0.8 0.8 0.8 
1 1 1 
0.09
0.032
873
1580
