0.300245 0.300245 0.514706 
0.2 0.2 0.2 
0.5 0.5 0.5 
1 1 1 
0.05 0.05 0.05 
0.8 0.8 0.8 
1 1 1 
0.09
0.032
1017
1920
