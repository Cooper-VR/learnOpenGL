0.0637255 0.0637255 0.0637255 
0 0 0 
0 0 0 
0 0 0 
0.102941 0.102941 0.102941 
1 1 1 
1 1 1 
0.09
0.032
0.05 0.05 0.05 
0.941176 0 0 
1 1 1 
0.09
0.032
0.808824 0.808824 0.808824 
0.8 0.8 0.8 
1 1 1 
0
0.032
0.05 0.05 0.05 
0.8 0.8 0.8 
1 1 1 
0.09
0.032
944
1702
